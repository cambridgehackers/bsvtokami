

`define HAZ BAZ
`HAZ;
`define N 2
typedef `N NUM_THINGS;

