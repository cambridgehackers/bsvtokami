import Vector::*, FIFO::*;
export Vector::*, FIFO::*;

// multiple variables
Bit#(32) a = 1, b = 2, c = 3;
