

module mkTest(Empty);
  Bit#(1) b = 22;
  let a = b;
endmodule