package BuildVector;

endpackage
