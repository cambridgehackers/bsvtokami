package StmtFSM;

endpackage
