package DefaultValue;

typeclass DefaultValue #( type t );
    t defaultValue ;
endtypeclass

endpackage
