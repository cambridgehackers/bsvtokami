package RevertingVirtualReg;

module mkRevertingVirtualReg#(a_type rst)(Reg#(a_type))
  provisos (Bits#(a_type, sizea));
endmodule

endpackage
