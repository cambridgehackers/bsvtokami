`define NumReadClients 1
`define NumWriteClients 1
`define PcieLanes 0
`define MemTagSize 12
`define SIM_DMA_READ_LATENCY 150
`define SIM_DMA_WRITE_LATENCY 150
`define TRACE_PORTAL 
`define ConnectalVersion 17.10.1
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 10
`define project_dir $(DTOP)
`define MainClockPeriod 8
`define DerivedClockPeriod 4.000000
`define PcieClockPeriod 8
`define XILINX 1
`define VirtexUltrascale 
`define PhysAddrWidth 40
`define DataBusWidth 128
`define XsimHostInterface 
`define AWSF1 1
`define DEFAULT_NOPROGRAM 1
`define CONNECTAL_BITS_DEPENDENCES build/checkpoints/to_aws/mkTop.SH_CL_routed.dcp
`define CONNECTAL_RUN_SCRIPT $(CONNECTALDIR)/scripts/run.aws
`define BOARD_awsf1 
