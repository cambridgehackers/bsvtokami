package Assert;
endpackage
