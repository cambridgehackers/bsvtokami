package Clocks;

interface Clock;
endinterface

interface Reset;
endinterface

module exposeCurrentClock(Clock);
endmodule

module exposeCurrentReset(Reset);
endmodule

endpackage
