typedef function a binop( a x, a y ) BinaryFunc#(type a);
