
import Foo::*;
import Foo::*;
import Foo::*, Baz::*;
export Foo::*;
export Bar(..);

export Baz::*, Fred(..);