
package FShow;
endpackage
