function Integer k(x,y)=3;
function Integer l(Integer x)=3;
module mkTest();
       function f();
        return ?;
       endfunction
       function g(Integer x);
        return ?;
       endfunction
       function h(x);
        return ?;
       endfunction
       function i;
        return ?;
       endfunction
       function Bool j;
        return ?;
       endfunction
       function d(x,y)=2;
       function Integer k(x,y)=3;
       function Integer l(Integer x)=3;
       function m provisos(Add#(1, 2, 3)) = 2;
endmodule


