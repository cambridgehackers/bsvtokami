

function Bool test_lt(Bit#(32) a, Bit#(32) b);
    return a < b;
endfunction
